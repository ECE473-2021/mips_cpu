// file forwarding_unit.v

module forwarding_unit(
	input wire ID_EX_RS,
	input wire ID_EX_RT,
	input wire EX_MEM_RD,
	input wire MEM_WB_RD,
	input wire EX_MEM_REGWRITE,
	input wire MEM_WB_REGWRITE,
	output reg ALU_A,
	output reg ALU_B
	);
	
	
endmodule
