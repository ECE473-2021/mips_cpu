// file forwarding_unit.v

module forwarding_unit(
	input wire ID_EX_RS,
	input wire ID_EX_RT,
	input wire EX_MEM_RD,
	input wire MEM_WB_RD,
	input wire EX_MEM_REGWRITE,
	input wire MEM_WB_REGWRITE,
	output wire ALU_A,
	output wire ALU_B
	);
	
	
endmodule
