// file ALU.v

module ALU(A,B,ALU_OP,ALU_OUT,ZERO);
	input wire [31:0] A,B;
	input wire [3:0] ALU_OP;
	output reg [31:0] ALU_OUT;
	output reg ZERO;
	
endmodule
